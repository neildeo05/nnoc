module ResultBuffer_int8 (clk, reset, result, res_buffer);

endmodule; // ResultBuffer_int8
